module core ();

    

endmodule //core