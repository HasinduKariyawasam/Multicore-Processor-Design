module ROM(addr,cs);

	input [4:0] addr;		// 5 bit address of microinstruction
	output [34:0] cs;		// Output 35-bit control signal
	
	reg [34:0] out;

	always @ (*)
		case (addr)
			5'd0: out = 35'b00001010000000000000000000000000001;	// FETCH1
			5'd1: out = 35'b010000000000000000000000000100xxxxx;	// FETCH2
			5'd2: out = 35'b00000000000000000000000000000100000;	// RSTALL1
			5'd3: out = 35'b00000010100001000000010111000000000;	// CONST1
			5'd4: out = 35'b10000000000000000000000000000000000;	// MOV1
			5'd5: out = 35'b00000100100001000000010111000000110;	// SIZE1
			5'd6: out = 35'b00000110000001000000010111000000111;	// SIZE2
			5'd7: out = 35'b00000011100001000000010111000001000;	// SIZE3
			5'd8: out = 35'b00000100000000000111010011000000000;	// SIZE4
			5'd9: out = 35'b00001010000000000000000000000001010;	// JMPNZY1
			5'd10: out = 35'b00000001101000000000000000000000000;	// JMPNZY2
			5'd11: out = 35'b00000000000000000000000000010000000;	// JMPNZN1
			5'd12: out = 35'b00000110000000001001001011000000000;	// MOV02_1
			5'd13: out = 35'b00000110000000001001001001000000000;	// MOV13_1
			5'd14: out = 35'b00000110000000100010100001000000000;	// ADDX1
			5'd15: out = 35'b00000110000000010010110001000000000;	// ADDY1
			5'd16: out = 35'b00000110000000000111010001000000000;	// ADD1
			5'd17: out = 35'b00000110000000000111010101000000000;	// SUB1
			5'd18: out = 35'b00000110000000000111010011000000000;	// MUL1
			5'd19: out = 35'b00000000111000000000000000000010100;	// LOAD1
			5'd20: out = 35'b00100001000000000000000000000000000;	// LOAD2
			5'd21: out = 35'b00000000111000000000000000000010110;	// STORE1
			5'd22: out = 35'b00000001010110000000000000000010111;	// STORE2
			5'd23: out = 35'b00010000000000000000000000000000000;	// STORE3
			5'd24: out = 35'b00000000000000000000000000100000000;	// INCI1
			5'd25: out = 35'b00000000000000000000000000001000000;	// RSTI1
			default: out = 35'd31; // Undefined microinstruction address - NOP
		endcase
	
	assign cs = out;
	
endmodule
