module ROM(addr,cs);

	input [4:0] addr;		// 5 bit address of microinstruction
	output [35:0] cs;		// Output 35-bit control signal
	
	reg [35:0] out;

	always @ (*)
		case (addr)
			5'd0: out = 36'b000010100000000000000000000000000001;	// FETCH1
			5'd1: out = 36'b0100000000000000000000000001000xxxxx;	// FETCH2
			5'd2: out = 36'b000000000000000000000000000001000000;	// RSTALL1
			5'd3: out = 36'b000000101000010000000101110000000000;	// CONST1
			5'd4: out = 36'b100000000000000000000000000000000000;	// MOV1
			5'd5: out = 36'b000001001000010000000101110000000110;	// SIZE1
			5'd6: out = 36'b000001100000010000000101110000000111;	// SIZE2
			5'd7: out = 36'b000000111000010000000101110000001000;	// SIZE3
			5'd8: out = 36'b000001000000000001110100010000000000;	// SIZE4
			5'd9: out = 36'b000010100000000000000000000000001010;	// JMPNZY1
			5'd10: out = 36'b000000011010000000000000000000000000;	// JMPNZY2
			5'd11: out = 36'b000000000000000000000000000100000000;	// JMPNZN1
			5'd12: out = 36'b000001100000000010010010110000000000;	// MOV02_1
			5'd13: out = 36'b000001100000000010010010010000000000;	// MOV13_1
			5'd14: out = 36'b000001100000001000101000010000000000;	// ADDX1
			5'd15: out = 36'b000001100000000100101100010000000000;	// ADDY1
			5'd16: out = 36'b000001100000000001110100010000000000;	// ADD1
			5'd17: out = 36'b000001100000000001110101010000000000;	// SUB1
			5'd18: out = 36'b000001100000000001110100110000000000;	// MUL1
			5'd19: out = 36'b000000001110000000000000000000010100;	// LOAD1
			5'd20: out = 36'b001000010000000000000000000000000000;	// LOAD2
			5'd21: out = 36'b000000001110000000000000000000010110;	// STORE1
			5'd22: out = 36'b000000010101100000000000000000010111;	// STORE2
			5'd23: out = 36'b000100000000000000000000000000000000;	// STORE3
			5'd24: out = 36'b000000000000000000000000001000000000;	// INCI1
			5'd25: out = 36'b000000000000000000000000000010000000;	// RSTI1
			5'd26: out = 36'b000000000000000000000000000000111111;	// OPEND1
			default: out = 36'd31; // Undefined microinstruction address - NOP
		endcase
	
	assign cs = out;
	
endmodule
