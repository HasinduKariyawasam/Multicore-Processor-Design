module ROM(addr,cs);

	input [4:0] addr;		// 5 bit address of microinstruction
	output [36:0] cs;		// 5 bit address of 1st microinstruction mapped from OPCODE address
	
	reg [36:0] out;

	always @ (*)
		case (addr)
			5'd0: out = 37'b0000001000000000000000000000000000001;	// FETCH1
			5'd1: out = 37'b01000100100000000000000000000100XXXXX;	// FETCH2
			5'd2: out = 37'b0000000000000000000000000000000100000;	// RSTALL1
			5'd3: out = 37'b0000000010100001000000010111000000000;	// CONST1
			5'd4: out = 37'b1000000000000000000000000000000000000;	// MOV1
			5'd5: out = 37'b0000000100100001000000010111000000110;	// SIZE1
			5'd6: out = 37'b0000000110000001000000010111000000111;	// SIZE2
			5'd7: out = 37'b0000000011100001000000010111000001000;	// SIZE3
			5'd8: out = 37'b0000000110000000000111010011000001001;	// SIZE4
			5'd9: out = 37'b0000000100011000000000000000000000000;	// SIZE5
			5'd10: out = 37'b0000001000000000000000000000000001011;	// JMPNZY1
			5'd11: out = 37'b0000010010000000000000000000010001100;	// JMPNZY2
			5'd12: out = 37'b0000000001101000000000000000000000000;	// JMPNZY3
			5'd13: out = 37'b0000000000000000000000000000010000000;	// JMPNZN1
			5'd14: out = 37'b0000000110000000001001001011000000000;	// MOVMSB1
			5'd15: out = 37'b0000000110000000001001001001000000000;	// MOVLSB1
			5'd16: out = 37'b0000000110000000100010100001000000000;	// ADDX1
			5'd17: out = 37'b0000000110000000010010110001000000000;	// ADDY1
			5'd18: out = 37'b0000000110000000000111010001000000000;	// ADD1
			5'd19: out = 37'b0000000110000000000111010101000000000;	// SUB1
			5'd20: out = 37'b0000000110000000000111010011000000000;	// MUL1
			5'd21: out = 37'b0001000000111000000000000000000010110;	// LOAD1
			5'd22: out = 37'b0010000001000000000000000000000000000;	// LOAD2
			5'd23: out = 37'b0000000000111000000000000000000011000;	// STORE1
			5'd24: out = 37'b0000100001010110000000000000000000000;	// STORE2
			5'd25: out = 37'b0000000000000000000000000000100000000;	// INCI1
			5'd26: out = 37'b0000000000000000000000000000001000000;	// RSTI1

		endcase
	
	assign cs = out;
	
endmodule
