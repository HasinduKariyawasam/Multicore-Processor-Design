module StoreController (input clk,
                        input opendFlag,
                        output memWrite, swEnable);
    
    wire regOut, startStore, storeEnd;

endmodule //StoreController